`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UCF KNIGHTS / NORTHROP GRUMMAN
// Engineer: Youssef Samwel
// Create Date: 11/19/2024 12:42:31 AM
//////////////////////////////////////////////////////////////////////////////////


module decoder_logic_testbench();



endmodule
