VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32b_1024_1rw_freepdk45
   CLASS BLOCK ;
   SIZE 237.8625 BY 216.5075 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  35.705 0.0 35.845 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.565 0.0 38.705 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.425 0.0 41.565 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.285 0.0 44.425 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.145 0.0 47.285 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.005 0.0 50.145 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.865 0.0 53.005 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  55.725 0.0 55.865 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.585 0.0 58.725 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.445 0.0 61.585 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.305 0.0 64.445 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.165 0.0 67.305 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.025 0.0 70.165 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  72.885 0.0 73.025 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  75.745 0.0 75.885 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.605 0.0 78.745 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.465 0.0 81.605 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.325 0.0 84.465 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.185 0.0 87.325 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.045 0.0 90.185 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  92.905 0.0 93.045 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  95.765 0.0 95.905 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  98.625 0.0 98.765 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.485 0.0 101.625 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.345 0.0 104.485 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.205 0.0 107.345 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.065 0.0 110.205 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  112.925 0.0 113.065 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  115.785 0.0 115.925 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  118.645 0.0 118.785 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  121.505 0.0 121.645 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  124.365 0.0 124.505 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.125 0.0 27.265 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  29.985 0.0 30.125 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  32.845 0.0 32.985 0.14 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 65.55 0.14 65.69 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 68.28 0.14 68.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 70.49 0.14 70.63 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 73.22 0.14 73.36 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 75.43 0.14 75.57 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 78.16 0.14 78.3 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 80.37 0.14 80.51 ;
      END
   END addr0[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 15.37 0.14 15.51 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 18.1 0.14 18.24 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 15.605 0.14 15.745 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  52.1075 0.0 52.2475 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.8275 0.0 57.9675 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  63.47 0.0 63.61 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  69.2675 0.0 69.4075 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.985 0.0 75.125 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.625 0.0 80.765 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  86.265 0.0 86.405 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  91.905 0.0 92.045 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  97.545 0.0 97.685 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  103.185 0.0 103.325 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.825 0.0 108.965 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.465 0.0 114.605 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.105 0.0 120.245 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  125.745 0.0 125.885 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.385 0.0 131.525 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  137.025 0.0 137.165 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  142.665 0.0 142.805 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  148.305 0.0 148.445 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  153.945 0.0 154.085 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  159.585 0.0 159.725 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  165.225 0.0 165.365 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  170.865 0.0 171.005 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  176.505 0.0 176.645 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  182.145 0.0 182.285 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  187.785 0.0 187.925 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  193.425 0.0 193.565 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.065 0.0 199.205 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  204.705 0.0 204.845 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  210.345 0.0 210.485 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.7225 23.0125 237.8625 23.1525 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.7225 22.5425 237.8625 22.6825 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.7225 22.7775 237.8625 22.9175 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  237.1625 0.0 237.8625 216.5075 ;
         LAYER metal3 ;
         RECT  0.0 0.0 237.8625 0.7 ;
         LAYER metal3 ;
         RECT  0.0 215.8075 237.8625 216.5075 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 216.5075 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 215.1075 ;
         LAYER metal3 ;
         RECT  1.4 1.4 236.4625 2.1 ;
         LAYER metal3 ;
         RECT  1.4 214.4075 236.4625 215.1075 ;
         LAYER metal4 ;
         RECT  235.7625 1.4 236.4625 215.1075 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 237.7225 216.3675 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 237.7225 216.3675 ;
   LAYER  metal3 ;
      RECT  0.28 65.41 237.7225 65.83 ;
      RECT  0.14 65.83 0.28 68.14 ;
      RECT  0.14 68.56 0.28 70.35 ;
      RECT  0.14 70.77 0.28 73.08 ;
      RECT  0.14 73.5 0.28 75.29 ;
      RECT  0.14 75.71 0.28 78.02 ;
      RECT  0.14 78.44 0.28 80.23 ;
      RECT  0.14 18.38 0.28 65.41 ;
      RECT  0.14 15.885 0.28 17.96 ;
      RECT  0.28 22.8725 237.5825 23.2925 ;
      RECT  0.28 23.2925 237.5825 65.41 ;
      RECT  237.5825 23.2925 237.7225 65.41 ;
      RECT  0.14 0.84 0.28 15.23 ;
      RECT  237.5825 0.84 237.7225 22.4025 ;
      RECT  0.14 80.65 0.28 215.6675 ;
      RECT  0.28 0.84 1.26 1.26 ;
      RECT  0.28 1.26 1.26 2.24 ;
      RECT  0.28 2.24 1.26 22.8725 ;
      RECT  1.26 0.84 236.6025 1.26 ;
      RECT  1.26 2.24 236.6025 22.8725 ;
      RECT  236.6025 0.84 237.5825 1.26 ;
      RECT  236.6025 1.26 237.5825 2.24 ;
      RECT  236.6025 2.24 237.5825 22.8725 ;
      RECT  0.28 65.83 1.26 214.2675 ;
      RECT  0.28 214.2675 1.26 215.2475 ;
      RECT  0.28 215.2475 1.26 215.6675 ;
      RECT  1.26 65.83 236.6025 214.2675 ;
      RECT  1.26 215.2475 236.6025 215.6675 ;
      RECT  236.6025 65.83 237.7225 214.2675 ;
      RECT  236.6025 214.2675 237.7225 215.2475 ;
      RECT  236.6025 215.2475 237.7225 215.6675 ;
   LAYER  metal4 ;
      RECT  35.425 0.42 36.125 216.3675 ;
      RECT  36.125 0.14 38.285 0.42 ;
      RECT  38.985 0.14 41.145 0.42 ;
      RECT  41.845 0.14 44.005 0.42 ;
      RECT  44.705 0.14 46.865 0.42 ;
      RECT  47.565 0.14 49.725 0.42 ;
      RECT  53.285 0.14 55.445 0.42 ;
      RECT  59.005 0.14 61.165 0.42 ;
      RECT  64.725 0.14 66.885 0.42 ;
      RECT  70.445 0.14 72.605 0.42 ;
      RECT  76.165 0.14 78.325 0.42 ;
      RECT  81.885 0.14 84.045 0.42 ;
      RECT  87.605 0.14 89.765 0.42 ;
      RECT  93.325 0.14 95.485 0.42 ;
      RECT  99.045 0.14 101.205 0.42 ;
      RECT  104.765 0.14 106.925 0.42 ;
      RECT  110.485 0.14 112.645 0.42 ;
      RECT  116.205 0.14 118.365 0.42 ;
      RECT  121.925 0.14 124.085 0.42 ;
      RECT  27.545 0.14 29.705 0.42 ;
      RECT  30.405 0.14 32.565 0.42 ;
      RECT  33.265 0.14 35.425 0.42 ;
      RECT  50.425 0.14 51.8275 0.42 ;
      RECT  52.5275 0.14 52.585 0.42 ;
      RECT  56.145 0.14 57.5475 0.42 ;
      RECT  58.2475 0.14 58.305 0.42 ;
      RECT  61.865 0.14 63.19 0.42 ;
      RECT  63.89 0.14 64.025 0.42 ;
      RECT  67.585 0.14 68.9875 0.42 ;
      RECT  69.6875 0.14 69.745 0.42 ;
      RECT  73.305 0.14 74.705 0.42 ;
      RECT  75.405 0.14 75.465 0.42 ;
      RECT  79.025 0.14 80.345 0.42 ;
      RECT  81.045 0.14 81.185 0.42 ;
      RECT  84.745 0.14 85.985 0.42 ;
      RECT  86.685 0.14 86.905 0.42 ;
      RECT  90.465 0.14 91.625 0.42 ;
      RECT  92.325 0.14 92.625 0.42 ;
      RECT  96.185 0.14 97.265 0.42 ;
      RECT  97.965 0.14 98.345 0.42 ;
      RECT  101.905 0.14 102.905 0.42 ;
      RECT  103.605 0.14 104.065 0.42 ;
      RECT  107.625 0.14 108.545 0.42 ;
      RECT  109.245 0.14 109.785 0.42 ;
      RECT  113.345 0.14 114.185 0.42 ;
      RECT  114.885 0.14 115.505 0.42 ;
      RECT  119.065 0.14 119.825 0.42 ;
      RECT  120.525 0.14 121.225 0.42 ;
      RECT  124.785 0.14 125.465 0.42 ;
      RECT  126.165 0.14 131.105 0.42 ;
      RECT  131.805 0.14 136.745 0.42 ;
      RECT  137.445 0.14 142.385 0.42 ;
      RECT  143.085 0.14 148.025 0.42 ;
      RECT  148.725 0.14 153.665 0.42 ;
      RECT  154.365 0.14 159.305 0.42 ;
      RECT  160.005 0.14 164.945 0.42 ;
      RECT  165.645 0.14 170.585 0.42 ;
      RECT  171.285 0.14 176.225 0.42 ;
      RECT  176.925 0.14 181.865 0.42 ;
      RECT  182.565 0.14 187.505 0.42 ;
      RECT  188.205 0.14 193.145 0.42 ;
      RECT  193.845 0.14 198.785 0.42 ;
      RECT  199.485 0.14 204.425 0.42 ;
      RECT  205.125 0.14 210.065 0.42 ;
      RECT  210.765 0.14 236.8825 0.42 ;
      RECT  0.98 0.14 26.845 0.42 ;
      RECT  0.98 0.42 1.12 1.12 ;
      RECT  0.98 1.12 1.12 215.3875 ;
      RECT  0.98 215.3875 1.12 216.3675 ;
      RECT  1.12 0.42 2.38 1.12 ;
      RECT  1.12 215.3875 2.38 216.3675 ;
      RECT  2.38 0.42 35.425 1.12 ;
      RECT  2.38 1.12 35.425 215.3875 ;
      RECT  2.38 215.3875 35.425 216.3675 ;
      RECT  36.125 0.42 235.4825 1.12 ;
      RECT  36.125 1.12 235.4825 215.3875 ;
      RECT  36.125 215.3875 235.4825 216.3675 ;
      RECT  235.4825 0.42 236.7425 1.12 ;
      RECT  235.4825 215.3875 236.7425 216.3675 ;
      RECT  236.7425 0.42 236.8825 1.12 ;
      RECT  236.7425 1.12 236.8825 215.3875 ;
      RECT  236.7425 215.3875 236.8825 216.3675 ;
   END
END    sram_32b_1024_1rw_freepdk45
END    LIBRARY
