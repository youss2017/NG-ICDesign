VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_150b_512_1rw_freepdk45
   CLASS BLOCK ;
   SIZE 485.975 BY 398.375 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.1075 0.0 54.2475 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.9675 0.0 57.1075 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.8275 0.0 59.9675 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.6875 0.0 62.8275 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.5475 0.0 65.6875 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.4075 0.0 68.5475 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.2675 0.0 71.4075 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.1275 0.0 74.2675 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.9875 0.0 77.1275 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.8475 0.0 79.9875 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.7075 0.0 82.8475 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.5675 0.0 85.7075 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.4275 0.0 88.5675 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  91.2875 0.0 91.4275 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  94.1475 0.0 94.2875 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  97.0075 0.0 97.1475 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.8675 0.0 100.0075 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.7275 0.0 102.8675 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  105.5875 0.0 105.7275 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.4475 0.0 108.5875 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  111.3075 0.0 111.4475 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.1675 0.0 114.3075 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  117.0275 0.0 117.1675 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.8875 0.0 120.0275 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  122.7475 0.0 122.8875 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  125.6075 0.0 125.7475 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  128.4675 0.0 128.6075 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.3275 0.0 131.4675 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  134.1875 0.0 134.3275 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  137.0475 0.0 137.1875 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  139.9075 0.0 140.0475 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  142.7675 0.0 142.9075 0.14 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  145.6275 0.0 145.7675 0.14 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  148.4875 0.0 148.6275 0.14 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  151.3475 0.0 151.4875 0.14 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  154.2075 0.0 154.3475 0.14 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  157.0675 0.0 157.2075 0.14 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  159.9275 0.0 160.0675 0.14 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  162.7875 0.0 162.9275 0.14 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  165.6475 0.0 165.7875 0.14 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  168.5075 0.0 168.6475 0.14 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  171.3675 0.0 171.5075 0.14 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  174.2275 0.0 174.3675 0.14 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  177.0875 0.0 177.2275 0.14 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  179.9475 0.0 180.0875 0.14 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  182.8075 0.0 182.9475 0.14 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  185.6675 0.0 185.8075 0.14 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  188.5275 0.0 188.6675 0.14 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.3875 0.0 191.5275 0.14 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  194.2475 0.0 194.3875 0.14 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.1075 0.0 197.2475 0.14 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.9675 0.0 200.1075 0.14 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  202.8275 0.0 202.9675 0.14 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  205.6875 0.0 205.8275 0.14 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  208.5475 0.0 208.6875 0.14 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.4075 0.0 211.5475 0.14 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  214.2675 0.0 214.4075 0.14 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  217.1275 0.0 217.2675 0.14 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  219.9875 0.0 220.1275 0.14 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  222.8475 0.0 222.9875 0.14 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  225.7075 0.0 225.8475 0.14 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.5675 0.0 228.7075 0.14 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  231.4275 0.0 231.5675 0.14 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  234.2875 0.0 234.4275 0.14 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  237.1475 0.0 237.2875 0.14 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  240.0075 0.0 240.1475 0.14 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  242.8675 0.0 243.0075 0.14 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  245.7275 0.0 245.8675 0.14 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  248.5875 0.0 248.7275 0.14 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  251.4475 0.0 251.5875 0.14 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  254.3075 0.0 254.4475 0.14 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  257.1675 0.0 257.3075 0.14 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.0275 0.0 260.1675 0.14 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  262.8875 0.0 263.0275 0.14 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  265.7475 0.0 265.8875 0.14 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  268.6075 0.0 268.7475 0.14 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  271.4675 0.0 271.6075 0.14 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  274.3275 0.0 274.4675 0.14 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  277.1875 0.0 277.3275 0.14 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  280.0475 0.0 280.1875 0.14 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  282.9075 0.0 283.0475 0.14 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  285.7675 0.0 285.9075 0.14 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  288.6275 0.0 288.7675 0.14 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  291.4875 0.0 291.6275 0.14 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  294.3475 0.0 294.4875 0.14 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  297.2075 0.0 297.3475 0.14 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  300.0675 0.0 300.2075 0.14 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  302.9275 0.0 303.0675 0.14 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  305.7875 0.0 305.9275 0.14 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  308.6475 0.0 308.7875 0.14 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  311.5075 0.0 311.6475 0.14 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  314.3675 0.0 314.5075 0.14 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  317.2275 0.0 317.3675 0.14 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  320.0875 0.0 320.2275 0.14 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  322.9475 0.0 323.0875 0.14 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  325.8075 0.0 325.9475 0.14 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  328.6675 0.0 328.8075 0.14 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  331.5275 0.0 331.6675 0.14 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  334.3875 0.0 334.5275 0.14 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  337.2475 0.0 337.3875 0.14 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  340.1075 0.0 340.2475 0.14 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  342.9675 0.0 343.1075 0.14 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  345.8275 0.0 345.9675 0.14 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  348.6875 0.0 348.8275 0.14 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  351.5475 0.0 351.6875 0.14 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  354.4075 0.0 354.5475 0.14 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  357.2675 0.0 357.4075 0.14 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  360.1275 0.0 360.2675 0.14 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  362.9875 0.0 363.1275 0.14 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  365.8475 0.0 365.9875 0.14 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  368.7075 0.0 368.8475 0.14 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  371.5675 0.0 371.7075 0.14 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  374.4275 0.0 374.5675 0.14 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  377.2875 0.0 377.4275 0.14 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  380.1475 0.0 380.2875 0.14 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  383.0075 0.0 383.1475 0.14 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  385.8675 0.0 386.0075 0.14 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  388.7275 0.0 388.8675 0.14 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  391.5875 0.0 391.7275 0.14 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  394.4475 0.0 394.5875 0.14 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  397.3075 0.0 397.4475 0.14 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  400.1675 0.0 400.3075 0.14 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  403.0275 0.0 403.1675 0.14 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  405.8875 0.0 406.0275 0.14 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  408.7475 0.0 408.8875 0.14 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  411.6075 0.0 411.7475 0.14 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  414.4675 0.0 414.6075 0.14 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  417.3275 0.0 417.4675 0.14 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  420.1875 0.0 420.3275 0.14 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  423.0475 0.0 423.1875 0.14 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  425.9075 0.0 426.0475 0.14 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  428.7675 0.0 428.9075 0.14 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  431.6275 0.0 431.7675 0.14 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  434.4875 0.0 434.6275 0.14 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  437.3475 0.0 437.4875 0.14 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  440.2075 0.0 440.3475 0.14 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  443.0675 0.0 443.2075 0.14 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  445.9275 0.0 446.0675 0.14 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  448.7875 0.0 448.9275 0.14 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  451.6475 0.0 451.7875 0.14 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  454.5075 0.0 454.6475 0.14 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  457.3675 0.0 457.5075 0.14 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  460.2275 0.0 460.3675 0.14 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  463.0875 0.0 463.2275 0.14 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  465.9475 0.0 466.0875 0.14 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  468.8075 0.0 468.9475 0.14 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  471.6675 0.0 471.8075 0.14 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  474.5275 0.0 474.6675 0.14 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  477.3875 0.0 477.5275 0.14 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  480.2475 0.0 480.3875 0.14 ;
      END
   END din0[149]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.2475 0.0 51.3875 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 78.02 0.14 78.16 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 80.75 0.14 80.89 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 82.96 0.14 83.1 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 85.69 0.14 85.83 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 87.9 0.14 88.04 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 90.63 0.14 90.77 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 92.84 0.14 92.98 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 95.57 0.14 95.71 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 22.38 0.14 22.52 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 25.11 0.14 25.25 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 22.615 0.14 22.755 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.09 0.0 79.23 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.8575 0.0 80.9975 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.95 0.0 82.09 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  83.6775 0.0 83.8175 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.81 0.0 84.95 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  86.4975 0.0 86.6375 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.67 0.0 87.81 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  89.3175 0.0 89.4575 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.4925 0.0 90.6325 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  92.1375 0.0 92.2775 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.3125 0.0 93.4525 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  94.9575 0.0 95.0975 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.25 0.0 96.39 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  97.7775 0.0 97.9175 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.11 0.0 99.25 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  100.5975 0.0 100.7375 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.97 0.0 102.11 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  103.4175 0.0 103.5575 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.8275 0.0 104.9675 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  106.2375 0.0 106.3775 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.6475 0.0 107.7875 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  109.0575 0.0 109.1975 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.4675 0.0 110.6075 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  111.8775 0.0 112.0175 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.2875 0.0 113.4275 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  114.6975 0.0 114.8375 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.1075 0.0 116.2475 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  117.5175 0.0 117.6575 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  118.9275 0.0 119.0675 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.3375 0.0 120.4775 0.14 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  121.7475 0.0 121.8875 0.14 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  123.1575 0.0 123.2975 0.14 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  124.5675 0.0 124.7075 0.14 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  125.9775 0.0 126.1175 0.14 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  127.3875 0.0 127.5275 0.14 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  128.7975 0.0 128.9375 0.14 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  130.2075 0.0 130.3475 0.14 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.6175 0.0 131.7575 0.14 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  133.0275 0.0 133.1675 0.14 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  134.4725 0.0 134.6125 0.14 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  135.8475 0.0 135.9875 0.14 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  137.3325 0.0 137.4725 0.14 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  138.6675 0.0 138.8075 0.14 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  140.1925 0.0 140.3325 0.14 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  141.4875 0.0 141.6275 0.14 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  143.0525 0.0 143.1925 0.14 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  144.3075 0.0 144.4475 0.14 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  145.9125 0.0 146.0525 0.14 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  147.1275 0.0 147.2675 0.14 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  148.7725 0.0 148.9125 0.14 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  149.9475 0.0 150.0875 0.14 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  151.6325 0.0 151.7725 0.14 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  152.7675 0.0 152.9075 0.14 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  154.4925 0.0 154.6325 0.14 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  155.5875 0.0 155.7275 0.14 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  157.3525 0.0 157.4925 0.14 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  158.4075 0.0 158.5475 0.14 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  160.39 0.0 160.53 0.14 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  161.2275 0.0 161.3675 0.14 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  163.21 0.0 163.35 0.14 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  164.0475 0.0 164.1875 0.14 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  164.89 0.0 165.03 0.14 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  166.8675 0.0 167.0075 0.14 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  167.75 0.0 167.89 0.14 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  169.6875 0.0 169.8275 0.14 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  170.61 0.0 170.75 0.14 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  172.5075 0.0 172.6475 0.14 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  173.47 0.0 173.61 0.14 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  175.3275 0.0 175.4675 0.14 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  176.33 0.0 176.47 0.14 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  178.1475 0.0 178.2875 0.14 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  179.19 0.0 179.33 0.14 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.9675 0.0 181.1075 0.14 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  182.05 0.0 182.19 0.14 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  183.7875 0.0 183.9275 0.14 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  184.91 0.0 185.05 0.14 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  186.6075 0.0 186.7475 0.14 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  187.77 0.0 187.91 0.14 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  189.4275 0.0 189.5675 0.14 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  190.6025 0.0 190.7425 0.14 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  192.2475 0.0 192.3875 0.14 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  193.4225 0.0 193.5625 0.14 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  195.0675 0.0 195.2075 0.14 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  196.35 0.0 196.49 0.14 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  197.8875 0.0 198.0275 0.14 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.21 0.0 199.35 0.14 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  200.7075 0.0 200.8475 0.14 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  202.07 0.0 202.21 0.14 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  203.5275 0.0 203.6675 0.14 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  204.93 0.0 205.07 0.14 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  206.3475 0.0 206.4875 0.14 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  207.7575 0.0 207.8975 0.14 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  209.1675 0.0 209.3075 0.14 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  210.5775 0.0 210.7175 0.14 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.9875 0.0 212.1275 0.14 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  213.3975 0.0 213.5375 0.14 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  214.8075 0.0 214.9475 0.14 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  216.2175 0.0 216.3575 0.14 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  217.6275 0.0 217.7675 0.14 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  219.0375 0.0 219.1775 0.14 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  220.4475 0.0 220.5875 0.14 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  221.8575 0.0 221.9975 0.14 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  223.2675 0.0 223.4075 0.14 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  224.6775 0.0 224.8175 0.14 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  226.0875 0.0 226.2275 0.14 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  227.4975 0.0 227.6375 0.14 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  228.9075 0.0 229.0475 0.14 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  230.3175 0.0 230.4575 0.14 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  231.7275 0.0 231.8675 0.14 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  233.1375 0.0 233.2775 0.14 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  234.5725 0.0 234.7125 0.14 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  235.9575 0.0 236.0975 0.14 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  237.44 0.0 237.58 0.14 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  238.7775 0.0 238.9175 0.14 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  240.2925 0.0 240.4325 0.14 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  241.5975 0.0 241.7375 0.14 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  243.1525 0.0 243.2925 0.14 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  244.4175 0.0 244.5575 0.14 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  246.0125 0.0 246.1525 0.14 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  247.2375 0.0 247.3775 0.14 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  248.8725 0.0 249.0125 0.14 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  250.0575 0.0 250.1975 0.14 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  251.7325 0.0 251.8725 0.14 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  252.8775 0.0 253.0175 0.14 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  254.5925 0.0 254.7325 0.14 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  255.6975 0.0 255.8375 0.14 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  257.4525 0.0 257.5925 0.14 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  258.5175 0.0 258.6575 0.14 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  260.5 0.0 260.64 0.14 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  261.3375 0.0 261.4775 0.14 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  263.32 0.0 263.46 0.14 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  264.1575 0.0 264.2975 0.14 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  266.14 0.0 266.28 0.14 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  266.9775 0.0 267.1175 0.14 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  267.85 0.0 267.99 0.14 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  269.7975 0.0 269.9375 0.14 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  270.71 0.0 270.85 0.14 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  272.6175 0.0 272.7575 0.14 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  273.57 0.0 273.71 0.14 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  275.4375 0.0 275.5775 0.14 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  276.43 0.0 276.57 0.14 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  278.2575 0.0 278.3975 0.14 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  279.29 0.0 279.43 0.14 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  281.0775 0.0 281.2175 0.14 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  282.15 0.0 282.29 0.14 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  283.8975 0.0 284.0375 0.14 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  285.01 0.0 285.15 0.14 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  286.7175 0.0 286.8575 0.14 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  287.87 0.0 288.01 0.14 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  289.5375 0.0 289.6775 0.14 ;
      END
   END dout0[149]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 398.375 ;
         LAYER metal3 ;
         RECT  0.0 397.675 485.975 398.375 ;
         LAYER metal3 ;
         RECT  0.0 0.0 485.975 0.7 ;
         LAYER metal4 ;
         RECT  485.275 0.0 485.975 398.375 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  483.875 1.4 484.575 396.975 ;
         LAYER metal3 ;
         RECT  1.4 396.275 484.575 396.975 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 396.975 ;
         LAYER metal3 ;
         RECT  1.4 1.4 484.575 2.1 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 485.835 398.235 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 485.835 398.235 ;
   LAYER  metal3 ;
      RECT  0.28 77.88 485.835 78.3 ;
      RECT  0.14 78.3 0.28 80.61 ;
      RECT  0.14 81.03 0.28 82.82 ;
      RECT  0.14 83.24 0.28 85.55 ;
      RECT  0.14 85.97 0.28 87.76 ;
      RECT  0.14 88.18 0.28 90.49 ;
      RECT  0.14 90.91 0.28 92.7 ;
      RECT  0.14 93.12 0.28 95.43 ;
      RECT  0.14 25.39 0.28 77.88 ;
      RECT  0.14 22.895 0.28 24.97 ;
      RECT  0.14 95.85 0.28 397.535 ;
      RECT  0.14 0.84 0.28 22.24 ;
      RECT  0.28 78.3 1.26 396.135 ;
      RECT  0.28 396.135 1.26 397.115 ;
      RECT  0.28 397.115 1.26 397.535 ;
      RECT  1.26 78.3 484.715 396.135 ;
      RECT  1.26 397.115 484.715 397.535 ;
      RECT  484.715 78.3 485.835 396.135 ;
      RECT  484.715 396.135 485.835 397.115 ;
      RECT  484.715 397.115 485.835 397.535 ;
      RECT  0.28 0.84 1.26 1.26 ;
      RECT  0.28 1.26 1.26 2.24 ;
      RECT  0.28 2.24 1.26 77.88 ;
      RECT  1.26 0.84 484.715 1.26 ;
      RECT  1.26 2.24 484.715 77.88 ;
      RECT  484.715 0.84 485.835 1.26 ;
      RECT  484.715 1.26 485.835 2.24 ;
      RECT  484.715 2.24 485.835 77.88 ;
   LAYER  metal4 ;
      RECT  53.8275 0.42 54.5275 398.235 ;
      RECT  54.5275 0.14 56.6875 0.42 ;
      RECT  57.3875 0.14 59.5475 0.42 ;
      RECT  60.2475 0.14 62.4075 0.42 ;
      RECT  63.1075 0.14 65.2675 0.42 ;
      RECT  65.9675 0.14 68.1275 0.42 ;
      RECT  68.8275 0.14 70.9875 0.42 ;
      RECT  71.6875 0.14 73.8475 0.42 ;
      RECT  74.5475 0.14 76.7075 0.42 ;
      RECT  291.9075 0.14 294.0675 0.42 ;
      RECT  294.7675 0.14 296.9275 0.42 ;
      RECT  297.6275 0.14 299.7875 0.42 ;
      RECT  300.4875 0.14 302.6475 0.42 ;
      RECT  303.3475 0.14 305.5075 0.42 ;
      RECT  306.2075 0.14 308.3675 0.42 ;
      RECT  309.0675 0.14 311.2275 0.42 ;
      RECT  311.9275 0.14 314.0875 0.42 ;
      RECT  314.7875 0.14 316.9475 0.42 ;
      RECT  317.6475 0.14 319.8075 0.42 ;
      RECT  320.5075 0.14 322.6675 0.42 ;
      RECT  323.3675 0.14 325.5275 0.42 ;
      RECT  326.2275 0.14 328.3875 0.42 ;
      RECT  329.0875 0.14 331.2475 0.42 ;
      RECT  331.9475 0.14 334.1075 0.42 ;
      RECT  334.8075 0.14 336.9675 0.42 ;
      RECT  337.6675 0.14 339.8275 0.42 ;
      RECT  340.5275 0.14 342.6875 0.42 ;
      RECT  343.3875 0.14 345.5475 0.42 ;
      RECT  346.2475 0.14 348.4075 0.42 ;
      RECT  349.1075 0.14 351.2675 0.42 ;
      RECT  351.9675 0.14 354.1275 0.42 ;
      RECT  354.8275 0.14 356.9875 0.42 ;
      RECT  357.6875 0.14 359.8475 0.42 ;
      RECT  360.5475 0.14 362.7075 0.42 ;
      RECT  363.4075 0.14 365.5675 0.42 ;
      RECT  366.2675 0.14 368.4275 0.42 ;
      RECT  369.1275 0.14 371.2875 0.42 ;
      RECT  371.9875 0.14 374.1475 0.42 ;
      RECT  374.8475 0.14 377.0075 0.42 ;
      RECT  377.7075 0.14 379.8675 0.42 ;
      RECT  380.5675 0.14 382.7275 0.42 ;
      RECT  383.4275 0.14 385.5875 0.42 ;
      RECT  386.2875 0.14 388.4475 0.42 ;
      RECT  389.1475 0.14 391.3075 0.42 ;
      RECT  392.0075 0.14 394.1675 0.42 ;
      RECT  394.8675 0.14 397.0275 0.42 ;
      RECT  397.7275 0.14 399.8875 0.42 ;
      RECT  400.5875 0.14 402.7475 0.42 ;
      RECT  403.4475 0.14 405.6075 0.42 ;
      RECT  406.3075 0.14 408.4675 0.42 ;
      RECT  409.1675 0.14 411.3275 0.42 ;
      RECT  412.0275 0.14 414.1875 0.42 ;
      RECT  414.8875 0.14 417.0475 0.42 ;
      RECT  417.7475 0.14 419.9075 0.42 ;
      RECT  420.6075 0.14 422.7675 0.42 ;
      RECT  423.4675 0.14 425.6275 0.42 ;
      RECT  426.3275 0.14 428.4875 0.42 ;
      RECT  429.1875 0.14 431.3475 0.42 ;
      RECT  432.0475 0.14 434.2075 0.42 ;
      RECT  434.9075 0.14 437.0675 0.42 ;
      RECT  437.7675 0.14 439.9275 0.42 ;
      RECT  440.6275 0.14 442.7875 0.42 ;
      RECT  443.4875 0.14 445.6475 0.42 ;
      RECT  446.3475 0.14 448.5075 0.42 ;
      RECT  449.2075 0.14 451.3675 0.42 ;
      RECT  452.0675 0.14 454.2275 0.42 ;
      RECT  454.9275 0.14 457.0875 0.42 ;
      RECT  457.7875 0.14 459.9475 0.42 ;
      RECT  460.6475 0.14 462.8075 0.42 ;
      RECT  463.5075 0.14 465.6675 0.42 ;
      RECT  466.3675 0.14 468.5275 0.42 ;
      RECT  469.2275 0.14 471.3875 0.42 ;
      RECT  472.0875 0.14 474.2475 0.42 ;
      RECT  474.9475 0.14 477.1075 0.42 ;
      RECT  477.8075 0.14 479.9675 0.42 ;
      RECT  51.6675 0.14 53.8275 0.42 ;
      RECT  77.4075 0.14 78.81 0.42 ;
      RECT  79.51 0.14 79.5675 0.42 ;
      RECT  80.2675 0.14 80.5775 0.42 ;
      RECT  81.2775 0.14 81.67 0.42 ;
      RECT  82.37 0.14 82.4275 0.42 ;
      RECT  83.1275 0.14 83.3975 0.42 ;
      RECT  84.0975 0.14 84.53 0.42 ;
      RECT  85.23 0.14 85.2875 0.42 ;
      RECT  85.9875 0.14 86.2175 0.42 ;
      RECT  86.9175 0.14 87.39 0.42 ;
      RECT  88.09 0.14 88.1475 0.42 ;
      RECT  88.8475 0.14 89.0375 0.42 ;
      RECT  89.7375 0.14 90.2125 0.42 ;
      RECT  90.9125 0.14 91.0075 0.42 ;
      RECT  91.7075 0.14 91.8575 0.42 ;
      RECT  92.5575 0.14 93.0325 0.42 ;
      RECT  93.7325 0.14 93.8675 0.42 ;
      RECT  94.5675 0.14 94.6775 0.42 ;
      RECT  95.3775 0.14 95.97 0.42 ;
      RECT  96.67 0.14 96.7275 0.42 ;
      RECT  97.4275 0.14 97.4975 0.42 ;
      RECT  98.1975 0.14 98.83 0.42 ;
      RECT  99.53 0.14 99.5875 0.42 ;
      RECT  100.2875 0.14 100.3175 0.42 ;
      RECT  101.0175 0.14 101.69 0.42 ;
      RECT  102.39 0.14 102.4475 0.42 ;
      RECT  103.8375 0.14 104.5475 0.42 ;
      RECT  105.2475 0.14 105.3075 0.42 ;
      RECT  106.6575 0.14 107.3675 0.42 ;
      RECT  108.0675 0.14 108.1675 0.42 ;
      RECT  109.4775 0.14 110.1875 0.42 ;
      RECT  110.8875 0.14 111.0275 0.42 ;
      RECT  112.2975 0.14 113.0075 0.42 ;
      RECT  113.7075 0.14 113.8875 0.42 ;
      RECT  115.1175 0.14 115.8275 0.42 ;
      RECT  116.5275 0.14 116.7475 0.42 ;
      RECT  117.9375 0.14 118.6475 0.42 ;
      RECT  119.3475 0.14 119.6075 0.42 ;
      RECT  120.7575 0.14 121.4675 0.42 ;
      RECT  122.1675 0.14 122.4675 0.42 ;
      RECT  123.5775 0.14 124.2875 0.42 ;
      RECT  124.9875 0.14 125.3275 0.42 ;
      RECT  126.3975 0.14 127.1075 0.42 ;
      RECT  127.8075 0.14 128.1875 0.42 ;
      RECT  129.2175 0.14 129.9275 0.42 ;
      RECT  130.6275 0.14 131.0475 0.42 ;
      RECT  132.0375 0.14 132.7475 0.42 ;
      RECT  133.4475 0.14 133.9075 0.42 ;
      RECT  134.8925 0.14 135.5675 0.42 ;
      RECT  136.2675 0.14 136.7675 0.42 ;
      RECT  137.7525 0.14 138.3875 0.42 ;
      RECT  139.0875 0.14 139.6275 0.42 ;
      RECT  140.6125 0.14 141.2075 0.42 ;
      RECT  141.9075 0.14 142.4875 0.42 ;
      RECT  143.4725 0.14 144.0275 0.42 ;
      RECT  144.7275 0.14 145.3475 0.42 ;
      RECT  146.3325 0.14 146.8475 0.42 ;
      RECT  147.5475 0.14 148.2075 0.42 ;
      RECT  149.1925 0.14 149.6675 0.42 ;
      RECT  150.3675 0.14 151.0675 0.42 ;
      RECT  152.0525 0.14 152.4875 0.42 ;
      RECT  153.1875 0.14 153.9275 0.42 ;
      RECT  154.9125 0.14 155.3075 0.42 ;
      RECT  156.0075 0.14 156.7875 0.42 ;
      RECT  157.7725 0.14 158.1275 0.42 ;
      RECT  158.8275 0.14 159.6475 0.42 ;
      RECT  160.81 0.14 160.9475 0.42 ;
      RECT  161.6475 0.14 162.5075 0.42 ;
      RECT  163.63 0.14 163.7675 0.42 ;
      RECT  164.4675 0.14 164.61 0.42 ;
      RECT  165.31 0.14 165.3675 0.42 ;
      RECT  166.0675 0.14 166.5875 0.42 ;
      RECT  167.2875 0.14 167.47 0.42 ;
      RECT  168.17 0.14 168.2275 0.42 ;
      RECT  168.9275 0.14 169.4075 0.42 ;
      RECT  170.1075 0.14 170.33 0.42 ;
      RECT  171.03 0.14 171.0875 0.42 ;
      RECT  171.7875 0.14 172.2275 0.42 ;
      RECT  172.9275 0.14 173.19 0.42 ;
      RECT  173.89 0.14 173.9475 0.42 ;
      RECT  174.6475 0.14 175.0475 0.42 ;
      RECT  175.7475 0.14 176.05 0.42 ;
      RECT  176.75 0.14 176.8075 0.42 ;
      RECT  177.5075 0.14 177.8675 0.42 ;
      RECT  178.5675 0.14 178.91 0.42 ;
      RECT  179.61 0.14 179.6675 0.42 ;
      RECT  180.3675 0.14 180.6875 0.42 ;
      RECT  181.3875 0.14 181.77 0.42 ;
      RECT  182.47 0.14 182.5275 0.42 ;
      RECT  183.2275 0.14 183.5075 0.42 ;
      RECT  184.2075 0.14 184.63 0.42 ;
      RECT  185.33 0.14 185.3875 0.42 ;
      RECT  186.0875 0.14 186.3275 0.42 ;
      RECT  187.0275 0.14 187.49 0.42 ;
      RECT  188.19 0.14 188.2475 0.42 ;
      RECT  188.9475 0.14 189.1475 0.42 ;
      RECT  189.8475 0.14 190.3225 0.42 ;
      RECT  191.0225 0.14 191.1075 0.42 ;
      RECT  191.8075 0.14 191.9675 0.42 ;
      RECT  192.6675 0.14 193.1425 0.42 ;
      RECT  193.8425 0.14 193.9675 0.42 ;
      RECT  194.6675 0.14 194.7875 0.42 ;
      RECT  195.4875 0.14 196.07 0.42 ;
      RECT  196.77 0.14 196.8275 0.42 ;
      RECT  197.5275 0.14 197.6075 0.42 ;
      RECT  198.3075 0.14 198.93 0.42 ;
      RECT  199.63 0.14 199.6875 0.42 ;
      RECT  200.3875 0.14 200.4275 0.42 ;
      RECT  201.1275 0.14 201.79 0.42 ;
      RECT  202.49 0.14 202.5475 0.42 ;
      RECT  203.9475 0.14 204.65 0.42 ;
      RECT  205.35 0.14 205.4075 0.42 ;
      RECT  206.7675 0.14 207.4775 0.42 ;
      RECT  208.1775 0.14 208.2675 0.42 ;
      RECT  209.5875 0.14 210.2975 0.42 ;
      RECT  210.9975 0.14 211.1275 0.42 ;
      RECT  212.4075 0.14 213.1175 0.42 ;
      RECT  213.8175 0.14 213.9875 0.42 ;
      RECT  215.2275 0.14 215.9375 0.42 ;
      RECT  216.6375 0.14 216.8475 0.42 ;
      RECT  218.0475 0.14 218.7575 0.42 ;
      RECT  219.4575 0.14 219.7075 0.42 ;
      RECT  220.8675 0.14 221.5775 0.42 ;
      RECT  222.2775 0.14 222.5675 0.42 ;
      RECT  223.6875 0.14 224.3975 0.42 ;
      RECT  225.0975 0.14 225.4275 0.42 ;
      RECT  226.5075 0.14 227.2175 0.42 ;
      RECT  227.9175 0.14 228.2875 0.42 ;
      RECT  229.3275 0.14 230.0375 0.42 ;
      RECT  230.7375 0.14 231.1475 0.42 ;
      RECT  232.1475 0.14 232.8575 0.42 ;
      RECT  233.5575 0.14 234.0075 0.42 ;
      RECT  234.9925 0.14 235.6775 0.42 ;
      RECT  236.3775 0.14 236.8675 0.42 ;
      RECT  237.86 0.14 238.4975 0.42 ;
      RECT  239.1975 0.14 239.7275 0.42 ;
      RECT  240.7125 0.14 241.3175 0.42 ;
      RECT  242.0175 0.14 242.5875 0.42 ;
      RECT  243.5725 0.14 244.1375 0.42 ;
      RECT  244.8375 0.14 245.4475 0.42 ;
      RECT  246.4325 0.14 246.9575 0.42 ;
      RECT  247.6575 0.14 248.3075 0.42 ;
      RECT  249.2925 0.14 249.7775 0.42 ;
      RECT  250.4775 0.14 251.1675 0.42 ;
      RECT  252.1525 0.14 252.5975 0.42 ;
      RECT  253.2975 0.14 254.0275 0.42 ;
      RECT  255.0125 0.14 255.4175 0.42 ;
      RECT  256.1175 0.14 256.8875 0.42 ;
      RECT  257.8725 0.14 258.2375 0.42 ;
      RECT  258.9375 0.14 259.7475 0.42 ;
      RECT  260.92 0.14 261.0575 0.42 ;
      RECT  261.7575 0.14 262.6075 0.42 ;
      RECT  263.74 0.14 263.8775 0.42 ;
      RECT  264.5775 0.14 265.4675 0.42 ;
      RECT  266.56 0.14 266.6975 0.42 ;
      RECT  267.3975 0.14 267.57 0.42 ;
      RECT  268.27 0.14 268.3275 0.42 ;
      RECT  269.0275 0.14 269.5175 0.42 ;
      RECT  270.2175 0.14 270.43 0.42 ;
      RECT  271.13 0.14 271.1875 0.42 ;
      RECT  271.8875 0.14 272.3375 0.42 ;
      RECT  273.0375 0.14 273.29 0.42 ;
      RECT  273.99 0.14 274.0475 0.42 ;
      RECT  274.7475 0.14 275.1575 0.42 ;
      RECT  275.8575 0.14 276.15 0.42 ;
      RECT  276.85 0.14 276.9075 0.42 ;
      RECT  277.6075 0.14 277.9775 0.42 ;
      RECT  278.6775 0.14 279.01 0.42 ;
      RECT  279.71 0.14 279.7675 0.42 ;
      RECT  280.4675 0.14 280.7975 0.42 ;
      RECT  281.4975 0.14 281.87 0.42 ;
      RECT  282.57 0.14 282.6275 0.42 ;
      RECT  283.3275 0.14 283.6175 0.42 ;
      RECT  284.3175 0.14 284.73 0.42 ;
      RECT  285.43 0.14 285.4875 0.42 ;
      RECT  286.1875 0.14 286.4375 0.42 ;
      RECT  287.1375 0.14 287.59 0.42 ;
      RECT  288.29 0.14 288.3475 0.42 ;
      RECT  289.0475 0.14 289.2575 0.42 ;
      RECT  289.9575 0.14 291.2075 0.42 ;
      RECT  0.98 0.14 50.9675 0.42 ;
      RECT  480.6675 0.14 484.995 0.42 ;
      RECT  54.5275 0.42 483.595 1.12 ;
      RECT  54.5275 1.12 483.595 397.255 ;
      RECT  54.5275 397.255 483.595 398.235 ;
      RECT  483.595 0.42 484.855 1.12 ;
      RECT  483.595 397.255 484.855 398.235 ;
      RECT  484.855 0.42 484.995 1.12 ;
      RECT  484.855 1.12 484.995 397.255 ;
      RECT  484.855 397.255 484.995 398.235 ;
      RECT  0.98 0.42 1.12 1.12 ;
      RECT  0.98 1.12 1.12 397.255 ;
      RECT  0.98 397.255 1.12 398.235 ;
      RECT  1.12 0.42 2.38 1.12 ;
      RECT  1.12 397.255 2.38 398.235 ;
      RECT  2.38 0.42 53.8275 1.12 ;
      RECT  2.38 1.12 53.8275 397.255 ;
      RECT  2.38 397.255 53.8275 398.235 ;
   END
END    sram_150b_512_1rw_freepdk45
END    LIBRARY
