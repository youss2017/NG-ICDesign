

module regfile (
    input  logic            i_clk,
    input  logic            i_reset,
    input  logic            i_rs1_out,
    input  logic            i_rs2_out,
    input  logic [4:0]      i_rs1,
    input  logic [4:0]      i_rs2, 
    input  logic [4:0]      i_rd,
    input  logic [31:0]     i_rd_data,
    output logic [XLEN-1:0] o_rs1_data,
    output logic [XLEN-1:0] o_rs2_data
);
    reg [XLEN-1:0] register_file [0:31];

    always_comb begin
        
        if (i_rs1_out) 
           if (i_rd == i_rs1)
               o_rs1_data = i_rd_data;
           else
               o_rs1_data = register_file[i_rs1];
        else 
            o_rs1_data = 'bz;
            
        if (i_rs2_out) 
           if (i_rd == i_rs2)
               o_rs2_data = i_rd_data;
           else
               o_rs2_data = register_file[i_rs2];
        else 
            o_rs2_data = 'bz;
                
    end

	always_ff @(posedge i_clk, posedge i_reset) begin
		if(i_reset) begin
            for(bit [4:0] i = 0; i < 32; i++)
                register_file[i] <= 0;
		end else begin
			if (i_rd > 0) 
				register_file[i_rd] <= i_rd_data;
		end
	end

endmodule