
// vcs -full64 -licqueue '-timescale=1ns/1ns' '+vcs+flush+all' '+warn=all' '-sverilog' \
//   '+incdir+%UVM_HOME%\src' %UVM_HOME%\src\uvm_pkg.sv -ntb_opts dtm -f files.f

// ./simv +vcs+lic+wait
// urg -dir simv.vdb -format both 
// ls -l urgReport\*.txt
// cat urgReport\*.txt
`timescale 1ns / 100ps

package rapid_pkg;

    parameter int XLEN = 32;

    parameter bit [XLEN-1:0] RESET_VECTOR = 0;
    parameter bit [XLEN-1:0] RESET_STACK_POINTER = 1024;
    parameter bit [XLEN-1:0] WORD_WIDTH = 4;
    parameter bit [XLEN-1:0] NOP_INSTRUCTION = 32'h00000033; // add x0, x0, x0
    parameter bit [XLEN-1:0] NOOP_INSTRUCTION = 32'h00000033; // add x0, x0, x0

    parameter bit [2:0] ADD_or_SUB = 3'b000;
    parameter bit [2:0] SLT = 3'b010;
    parameter bit [2:0] SLTU = 3'b011;
    parameter bit [2:0] XOR_ = 3'b100;
    parameter bit [2:0] OR_ = 3'b110;
    parameter bit [2:0] AND_ = 3'b111;
    parameter bit [2:0] SLL = 3'b001;
    parameter bit [2:0] SRL_or_SRA = 3'b101;
    parameter bit [2:0] LB_or_SB = 3'b000;
    parameter bit [2:0] LH_or_SH = 3'b001;
    parameter bit [2:0] LW_or_SW = 3'b010;
    parameter bit [2:0] LBU = 3'b100;
    parameter bit [2:0] LHU = 3'b101;
    parameter bit [2:0] BLTU = 3'b110;
    parameter bit [2:0] BGEU = 3'b111;

    // this is the largest control signal
    // its generated by the decoder and used by
    // the execute stage.
    typedef struct {
        logic load_upper_imm;
        logic uncond_branch;
        logic cond_branch;
        logic mem;
        logic alu_imm;
        logic alu_reg;
        logic iop;
        logic rs1_out;
        logic rs2_out;
        logic [2:0] fcs_opcode;
        logic [4:0] rs1;
        logic [4:0] rs2;
        logic [4:0] rd;
        logic [XLEN-1:0] debug_instruction;
    } control_ex_s;

    // Control signal for cpu memory stage
    typedef struct {
        logic mem;
        logic iop;
        logic [2:0] fcs_opcode;
        logic [4:0] rd;
        logic [XLEN-1:0] debug_instruction;
    } control_mem_s;
    

    // Define a default state function for control_s
    function automatic control_ex_s control_ex_s_default();
        control_ex_s_default = '{ 
            load_upper_imm: '0,
            uncond_branch: '0,
            cond_branch: '0,
            mem: '0,
            alu_imm: '0,
            alu_reg: '0,
            iop: '0,
            rs1_out: '0,
            rs2_out: '0,
            fcs_opcode: '0,
            rs1: '0,
            rs2: '0,
            rd: '0,
            debug_instruction: 'x
        };
    endfunction

        // Define a default state function for control_s
    function automatic control_mem_s control_mem_s_default();
        control_mem_s_default = '{ 
            mem: '0,
            iop: '0,
            fcs_opcode: '0,
            rd: '0,
            debug_instruction: 'x
        };
    endfunction

    
endpackage

import rapid_pkg::*;

module execute_state

(
    input logic                          i_clk,
    input logic                          i_reset,
    input logic                          i_pc_load,
    input logic         [XLEN-1:0]       i_pc,
    input control_ex_s                   i_control_signal,
    input logic signed  [XLEN-1:0]       i_rs1,
    input logic signed  [XLEN-1:0]       i_rs2,
    input logic signed  [XLEN-1:0]       i_imm,
    output logic        [XLEN-1:0]       o_pc,
    output control_ex_s                  o_control_signal,
    output logic signed  [XLEN-1:0]      o_rs1,
    output logic signed  [XLEN-1:0]      o_rs2,
  output logic signed  [XLEN-1:0]      o_imm
);

    // internal value
    control_ex_s iv_control_signal;
    logic signed [XLEN-1:0] iv_rs1, iv_rs2, iv_imm, iv_pc;

    assign o_pc             = iv_pc;
    assign o_control_signal = iv_control_signal;
    assign o_rs1            = iv_rs1;
    assign o_rs2            = iv_rs2;
    assign o_imm            = iv_imm;

    always_ff @(posedge i_clk, posedge i_reset) begin

        if (i_reset) begin
            iv_control_signal <= control_ex_s_default();
            iv_rs1            <= 0;
            iv_rs2            <= 0;
            iv_imm            <= 0;
            iv_pc             <= 0;
        end else begin
            // Load data from inputs ports to local state
            iv_pc               <= i_pc_load ?  0                       : i_pc;
            iv_control_signal   <= i_pc_load ?  control_ex_s_default()  : i_control_signal;
            iv_rs1              <= i_pc_load ?  0                       : i_rs1;
            iv_rs2              <= i_pc_load ?  0                       : i_rs2;
            iv_imm              <= i_pc_load ?  0                       : i_imm;
        end        

    end


endmodule

import rapid_pkg::*;

module execute_logic
(
    input  logic                       i_clk,
    input  logic        [XLEN-1:0]     i_pc,
    input  control_ex_s                i_control_signal,
    input  logic signed [XLEN-1:0]     i_rs1,
    input  logic signed [XLEN-1:0]     i_rs2,
    input  logic signed [XLEN-1:0]     i_imm,
    output control_mem_s               o_control_signal,
    output logic                       o_pc_load,
    output logic        [XLEN-1:0]     o_pc_ext,
    output logic        [XLEN-1:0]     o_memory_data,
    output logic        [XLEN-1:0]     o_rd_output
);

    // We’ll store the outputs in internal registers (or logic variables).
    // Then we assign them to the module outputs at the bottom.
    control_mem_s r_control_signal;
    logic         r_pc_load;
    logic [XLEN-1:0] r_pc_ext;
    logic [XLEN-1:0] r_memory_data;
  logic [XLEN-1:0] r_rd_output;

    // "Wire" for the second ALU operand selection
    wire [XLEN-1:0] port2 = (i_control_signal.alu_reg) ? i_rs2 : i_imm;

    // Assign output ports from internal registers
    assign o_control_signal = r_control_signal;
    assign o_pc_load        = r_pc_load;
    assign o_pc_ext         = r_pc_ext;
    assign o_memory_data    = r_memory_data;
    assign o_rd_output      = r_rd_output;


    // Sequential: Update outputs on rising clock edge
    always_ff @(posedge i_clk) begin

        // Default assignments each clock
        r_control_signal.mem              <= i_control_signal.mem;
        r_control_signal.iop              <= i_control_signal.iop;
        r_control_signal.fcs_opcode       <= i_control_signal.fcs_opcode;
        r_control_signal.rd               <= i_control_signal.rd;
        r_control_signal.debug_instruction<= i_control_signal.debug_instruction;

        r_pc_load  <= 1'b0;
        r_pc_ext   <= 0;
        r_rd_output <= 0;

        // For convenience, memory_data is always the i_rs2 value
        r_memory_data <= i_rs2;

        // ALU (Register or Immediate)
        if (i_control_signal.alu_imm || i_control_signal.alu_reg) begin
            case (i_control_signal.fcs_opcode)
                ADD_or_SUB: r_rd_output <= (i_control_signal.iop) 
                                         ? (i_rs1 - port2) 
                                         : (i_rs1 + port2);
                SLT:        r_rd_output <= (i_rs1 < port2) ? 1 : 0;
                SLTU:       r_rd_output <= ($unsigned(i_rs1) < $unsigned(port2)) ? 1 : 0;
                XOR_:       r_rd_output <= i_rs1 ^ port2;
                OR_:        r_rd_output <= i_rs1 | port2;
                AND_:       r_rd_output <= i_rs1 & port2;
                SLL:        r_rd_output <= i_rs1 << port2[4:0];
                SRL_or_SRA: begin
                                if (!i_control_signal.iop)
                                    r_rd_output <= i_rs1 >> port2[4:0];
                                else
                                    r_rd_output <= i_rs1 >>> port2[4:0];
                            end
                default:    r_rd_output <= 0; 
            endcase

            // No PC update in an ALU instruction
            r_pc_load <= 1'b0;
            r_pc_ext  <= 0;
        end

      // Conditional Branch
        else if (i_control_signal.cond_branch) begin
            case (i_control_signal.fcs_opcode)
                3'b000 /*BEQ*/:  r_pc_load <= (i_rs1 == i_rs2);
                3'b001 /*BNE*/:  r_pc_load <= (i_rs1 != i_rs2);
                3'b100 /*BLT*/:  r_pc_load <= (i_rs1 <  i_rs2);
                3'b101 /*BGE*/:  r_pc_load <= (i_rs1 >= i_rs2);
                3'b110 /*BLTU*/: r_pc_load <= ($unsigned(i_rs1) <  $unsigned(i_rs2));
                3'b111 /*BGEU*/: r_pc_load <= ($unsigned(i_rs1) >= $unsigned(i_rs2));
                default:         r_pc_load <= 1'b0;
            endcase
            r_pc_ext  <= (i_pc + i_imm) & ~32'h1;
        end

        // Unconditional Branch
        else if (i_control_signal.uncond_branch) begin
            // rd gets PC+4
            r_rd_output <= i_pc + 4;
            // JALR vs. JAL
            if (i_control_signal.iop)
                r_pc_ext <= (i_rs1 + i_imm) & ~32'h1;  // JALR
            else
                r_pc_ext <= (i_pc + i_imm)  & ~32'h1;  // JAL
            r_pc_load <= 1'b1;
        end

        // LUI & AUIPC
        else if (i_control_signal.load_upper_imm) begin
            if (i_control_signal.iop) 
                // LUI
                r_rd_output <= i_imm;
            else 
                // AUIPC
                r_rd_output <= i_pc + i_imm;
            r_pc_ext  <= 0;
            r_pc_load <= 1'b0;
        end

        // Memory Operations
        else if (i_control_signal.mem) begin
            r_rd_output <= i_rs1 + i_imm;
            r_pc_ext    <= 0;
            r_pc_load   <= 1'b0;
        end

        // Default / NOP
        else begin
            r_pc_load   <= 1'b0;
            r_pc_ext    <= 0;
            r_rd_output <= 0;
        end
    end

endmodule